/*
Reacts to drift events - Allows drifts to offset the next limit during preemptive events. 
Uses active High Half-Rate and Low Half-Rate during event updates.
*/