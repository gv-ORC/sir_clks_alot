package common_p;

    typedef struct packed {
        logic clk;
        logic clk_en;
        logic sync_rst;
    } clk_dom_s;

endpackage
